module logic(input wire[15:0] in_a, input wire[15:0] in_b, input wire[3:0] sel);
	always_comb begin
		case(sel)
			
		endcase
	end
endmodule
