interface alu_if (
    input logic clk
);

  //input_1
  logic [15:0] in_a;
  //input_2
  logic [15:0] in_b;
  //output
  logic [15:0] out;
endinterface
