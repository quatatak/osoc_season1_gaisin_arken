module top_module(input wire carry_in, input wire[15:0] in_a, input wire[15:0] in_b, input wire[3:0] select, input wire mode, output wire[15:0] alu_out, output wire carry_out, output wire compare);
	
endmodule
