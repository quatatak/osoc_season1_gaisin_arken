typedef uvm_sequencer#(alu_packet) alu_sequencer;

